`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    10:24:28 09/01/2014 
// Design Name: 
// Module Name:    Masking_Module 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module Masking_Module(
input[63:0] A,
input[7:0] B,
output  [63:0] Out

    );
assign Out=(B==8'h1)?({A[63:1],1'h0}):
           ((B==8'h2)?({A[63:2],2'h0}):
           ((B==8'h3)?({A[63:3],3'h0}):
           ((B==8'h4)?({A[63:4],4'h0}):
           ((B==8'h5)?({A[63:5],5'h0}):
           ((B==8'h6)?({A[63:6],6'h0}):
           ((B==8'h7)?({A[63:7],7'h0}):
           ((B==8'h8)?({A[63:8],8'h0}):	
            ((B==8'h9)?({A[63:9],9'h0}):
           ((B==8'ha)?({A[63:10],10'h0}):
           ((B==8'hb)?({A[63:11],11'h0}):
           ((B==8'hc)?({A[63:12],12'h0}):
           ((B==8'hd)?({A[63:13],13'h0}):
           ((B==8'he)?({A[63:14],14'h0}):
           ((B==8'hf)?({A[63:15],15'h0}):	
            ((B==8'h10)?({A[63:16],16'h0}):
           ((B==8'h11)?({A[63:17],17'h0}):
           ((B==8'h12)?({A[63:18],18'h0}):
           ((B==8'h13)?({A[63:19],19'h0}):
           ((B==8'h14)?({A[63:20],20'h0}):
           ((B==8'h15)?({A[63:21],21'h0}):
           ((B==8'h16)?({A[63:22],22'h0}):
            ((B==8'h17)?({A[63:23],23'h0}):
           ((B==8'h18)?({A[63:24],24'h0}):
           ((B==8'h19)?({A[63:25],25'h0}):
           ((B==8'h1a)?({A[63:26],26'h0}):
           ((B==8'h1b)?({A[63:27],27'h0}):
           ((B==8'h1c)?({A[63:28],28'h0}):
           ((B==8'h1d)?({A[63:29],29'h0}):	
			  ((B==8'h1e)?({A[63:30],30'h0}):
           ((B==8'h1f)?({A[63:31],31'h0}):
           ((B==8'h20)?({A[63:32],32'h0}):
           ((B==8'h21)?({A[63:33],33'h0}):
           ((B==8'h22)?({A[63:34],34'h0}):
           ((B==8'h23)?({A[63:35],35'h0}):
           ((B==8'h24)?({A[63:36],36'h0}):	
           ((B==8'h25)?({A[63:37],37'h0}):
           ((B==8'h26)?({A[63:38],38'h0}):
           ((B==8'h27)?({A[63:39],39'h0}):
           ((B==8'h28)?({A[63:40],40'h0}):
           ((B==8'h29)?({A[63:41],41'h0}):
           ((B==8'h2a)?({A[63:42],42'h0}):
           ((B==8'h2b)?({A[63:43],43'h0}):	
           ((B==8'h2c)?({A[63:44],44'h0}):
           ((B==8'h2d)?({A[63:45],45'h0}):
           ((B==8'h2e)?({A[63:46],46'h0}):
           ((B==8'h2f)?({A[63:47],47'h0}):
           ((B==8'h30)?({A[63:48],48'h0}):
           ((B==8'h31)?({A[63:49],49'h0}):
           ((B==8'h32)?({A[63:50],50'h0}):
           ((B==8'h33)?({A[63:51],51'h0}):
           ((B==8'h34)?({A[63:52],52'h0}):
           ((B==8'h35)?({A[63:53],53'h0}):
           ((B==8'h36)?({A[63:54],54'h0}):
           ((B==8'h37)?({A[63:55],55'h0}):
           ((B==8'h38)?({A[63:56],56'h0}):
           ((B==8'h39)?({A[63:57],57'h0}):	
			  ((B==8'h3a)?({A[63:58],58'h0}):
           ((B==8'h3b)?({A[63:59],59'h0}):
           ((B==8'h3c)?({A[63:60],60'h0}):
           ((B==8'h3d)?({A[63:61],61'h0}):
           ((B==8'h3e)?({A[63:62],62'h0}):
           ((B==8'h3f)?({A[63],63'h0}):A))))))))))))))))))))))))))))))))))))))))))))))))))))))))))))));
           			  
endmodule
